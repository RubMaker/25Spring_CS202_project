`timescale 1ns / 1ps
`include "Constants.vh"



module VGADisplay (
    input wire clk,
    input wire reset_n,

    //input wire [7:0] script, // 8switch
    
    input wire [7:0] data, // datain
    //input wire [7:0] led_2, // 8led_right

    
    /*input wire [7:0] segment0,
    input wire [7:0] segment1,
    input wire [7:0] segment2,
    input wire [7:0] segment3,
    input wire [7:0] segment4,
    input wire [7:0] segment5,
    input wire [7:0] segment6,
    input wire [7:0] segment7,*/

    
    
    //input wire [7:0] game_mode, //state
    output hsync,   // line synchronization signal
    output vsync,   // vertical synchronization signal
    output reg [3:0] red,
    output reg [3:0] green,
    output reg [3:0] blue
);

//num_none: nothing
//num_zero-num_nine: 32x32 pixel font for numbers 0-9
//char_dai:��
//char_ding:��
//char_mo:ģ
//char_shi:ʽ
//char_ji:��
//char_suan:��
//char_xue:ѧ
//char_xi:ϰ
//char_yan:��
//char_shi2:ʾ
//char_dui:��
//char_cuo:��
//char_guan:��
//char_ji2:��

/*parameter [0:1023] char_none={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};*/
parameter [0:1023] num_zero={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00111110, 8'b00001111, 8'b10000000, 8'b00000000, 
    8'b00111100, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00111110, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00111111, 8'b00001111, 8'b10000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};

parameter [0:1023] num_one={
     8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b01111111, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b01111111, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b01111011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b01100011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};/*

parameter [0:1023] num_two={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00111110, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00111110, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111000, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00001111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00011111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00111111, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11100000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b10000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111110, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b01111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b01111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};

parameter [0:1023] num_three={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00111110, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00001111, 8'b10000000, 8'b00000000, 
    8'b00000001, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00000001, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111110, 8'b00001111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};

parameter [0:1023] num_four={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00011110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00111110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b01111110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11101110, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11001110, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b10001110, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b10001110, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b00111110, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b01111100, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b11111000, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b11111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b11111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b11111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00000000, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};

parameter num_five={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111101, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00111110, 8'b00001111, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111110, 8'b00001111, 8'b10000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};

parameter [0:1023] num_six={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00011111, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00111110, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b01111000, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b01111011, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b01111111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b01111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b01111111, 8'b00001111, 8'b11000000, 8'b00000000, 
    8'b01111110, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b00001111, 8'b10000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00001111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};

parameter [0:1023] num_seven={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b11111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b11111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b11111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b11111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00001111, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00001111, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00011111, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00011110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00111110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00111100, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00111100, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b01111100, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b11110000, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11110000, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11110000, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11100000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11100000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b10000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};

parameter [0:1023] num_eight={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b10111111, 8'b10000000, 8'b00000000, 
    8'b00111110, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b01111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111110, 8'b00001111, 8'b10000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00001111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b01111110, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11100000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11100000, 8'b00000000, 
    8'b01111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111110, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00001111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};

parameter [0:1023] num_nine={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00111110, 8'b00001111, 8'b10000000, 8'b00000000, 
    8'b01111100, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b01111000, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b00011111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00000111, 8'b11111011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b11000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00111100, 8'b00001111, 8'b10000000, 8'b00000000, 
    8'b00111110, 8'b00011111, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11110000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};

parameter [0:1023] char_neg={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b01111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b01111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b01111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};
parameter [0:1023] char_A={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11011110, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11011111, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11011111, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b10001111, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b10001111, 8'b10000000, 8'b00000000, 
    8'b00001111, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00001111, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00011111, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00011110, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b01111100, 8'b00000001, 8'b11110000, 8'b00000000, 
    8'b01111000, 8'b00000000, 8'b11110000, 8'b00000000, 
    8'b11111000, 8'b00000000, 8'b11111000, 8'b00000000, 
    8'b11111000, 8'b00000000, 8'b11111000, 8'b00000000, 
    8'b11110000, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b11110000, 8'b00000000, 8'b01111100, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};
parameter [0:1023] char_B={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11110000, 8'b00000000, 
    8'b00111100, 8'b00000001, 8'b11110000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b11110000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b11110000, 8'b00000000, 
    8'b00111100, 8'b00000001, 8'b11110000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11110000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11110000, 8'b00000000, 
    8'b00111100, 8'b00000001, 8'b11111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b11111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b11111000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11111000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11110000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};
parameter [0:1023] char_C={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00000011, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00001111, 8'b11111111, 8'b11110000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b11111000, 8'b00000000, 
    8'b00011111, 8'b10000001, 8'b11111000, 8'b00000000, 
    8'b00111111, 8'b00000000, 8'b01111100, 8'b00000000, 
    8'b00111110, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b01111100, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b01111100, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b01111000, 8'b00000000, 8'b00011100, 8'b00000000, 
    8'b01111100, 8'b00000000, 8'b00111110, 8'b00000000, 
    8'b01111100, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b00111110, 8'b00000000, 8'b01111100, 8'b00000000, 
    8'b00111111, 8'b00000000, 8'b11111100, 8'b00000000, 
    8'b00011111, 8'b10000001, 8'b11111000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b11110000, 8'b00000000, 
    8'b00001111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00000011, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};
parameter [0:1023] char_D={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11110000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111100, 8'b00000111, 8'b11110000, 8'b00000000, 
    8'b00111100, 8'b00000001, 8'b11110000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b11111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b01111100, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b11111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b11111000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11110000, 8'b00000000, 
    8'b00111100, 8'b00001111, 8'b11110000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};
parameter [0:1023] char_E={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11110000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11110000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11110000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};
parameter [0:1023] char_F={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};
parameter [0:1023] char_guan={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b01100000, 8'b00000111, 8'b10000000, 
    8'b00000001, 8'b11100000, 8'b00000111, 8'b10000000, 
    8'b00000001, 8'b11110000, 8'b00001111, 8'b00000000, 
    8'b00000000, 8'b11111000, 8'b00001111, 8'b00000000, 
    8'b00000000, 8'b01111000, 8'b00011111, 8'b00000000, 
    8'b00000000, 8'b01111100, 8'b00011110, 8'b00000000, 
    8'b00000000, 8'b00111100, 8'b00111110, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00000000, 8'b00001111, 8'b11100000, 8'b00000000, 
    8'b00000000, 8'b00001111, 8'b11110000, 8'b00000000, 
    8'b00000000, 8'b00011111, 8'b11111000, 8'b00000000, 
    8'b00000000, 8'b00011110, 8'b01111100, 8'b00000000, 
    8'b00000000, 8'b00111110, 8'b01111110, 8'b00000000, 
    8'b00000000, 8'b01111100, 8'b00111111, 8'b00000000, 
    8'b00000001, 8'b11111100, 8'b00011111, 8'b10000000, 
    8'b00000111, 8'b11110000, 8'b00001111, 8'b11100000, 
    8'b00011111, 8'b11100000, 8'b00000111, 8'b11111100, 
    8'b01111111, 8'b11000000, 8'b00000001, 8'b11111110, 
    8'b01111111, 8'b00000000, 8'b00000000, 8'b11111110, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00111100, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00001100
};

parameter [0:1023] char_ji2={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000001, 8'b11111111, 8'b11000000, 
    8'b00000011, 8'b11000011, 8'b11111111, 8'b11000000, 
    8'b00000011, 8'b11000011, 8'b11111111, 8'b11000000, 
    8'b00000011, 8'b11000011, 8'b11111111, 8'b11000000, 
    8'b00000011, 8'b11000011, 8'b11000011, 8'b11000000, 
    8'b01111111, 8'b11111111, 8'b11000011, 8'b11000000, 
    8'b01111111, 8'b11111111, 8'b11000011, 8'b11000000, 
    8'b01111111, 8'b11111111, 8'b11000011, 8'b11000000, 
    8'b01111111, 8'b11111111, 8'b11000011, 8'b11000000, 
    8'b00000111, 8'b11000011, 8'b11000011, 8'b11000000, 
    8'b00000111, 8'b11100011, 8'b11000011, 8'b11000000, 
    8'b00001111, 8'b11110011, 8'b11000011, 8'b11000000, 
    8'b00001111, 8'b11111011, 8'b11000011, 8'b11000000, 
    8'b00001111, 8'b11111011, 8'b11000011, 8'b11000000, 
    8'b00011111, 8'b11111111, 8'b11000011, 8'b11000000, 
    8'b00111111, 8'b11111111, 8'b11000011, 8'b11000000, 
    8'b00111111, 8'b11011011, 8'b11000011, 8'b11000000, 
    8'b01111011, 8'b11011011, 8'b11000011, 8'b11000000, 
    8'b01111011, 8'b11000011, 8'b11000011, 8'b11000000, 
    8'b01110011, 8'b11000011, 8'b11000011, 8'b11001110, 
    8'b01110011, 8'b11000011, 8'b10000011, 8'b11001110, 
    8'b01100011, 8'b11000111, 8'b10000011, 8'b11001110, 
    8'b00000011, 8'b11000111, 8'b10000011, 8'b11001110, 
    8'b00000011, 8'b11000111, 8'b10000011, 8'b11001110, 
    8'b00000011, 8'b11001111, 8'b00000011, 8'b11001110, 
    8'b00000011, 8'b11011111, 8'b00000011, 8'b11111110, 
    8'b00000011, 8'b11011111, 8'b00000011, 8'b11111110, 
    8'b00000011, 8'b11011110, 8'b00000001, 8'b11111110, 
    8'b00000011, 8'b11011110, 8'b00000000, 8'b11111100, 
    8'b00000011, 8'b10001100, 8'b00000000, 8'b00000000
};

parameter [0:1023] char_dai={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11000000, 8'b00011110, 8'b00000000, 
    8'b00000011, 8'b11100000, 8'b00011110, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b11001111, 8'b11111111, 8'b11111100, 
    8'b00001111, 8'b10001111, 8'b11111111, 8'b11111100, 
    8'b00011111, 8'b00001111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b00001111, 8'b11111111, 8'b11111100, 
    8'b01111110, 8'b11000000, 8'b00011110, 8'b00000000, 
    8'b01111100, 8'b11110000, 8'b00011110, 8'b00000000, 
    8'b01111001, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b01110011, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00000011, 8'b11011111, 8'b11111111, 8'b11111110, 
    8'b00000111, 8'b11011111, 8'b11111111, 8'b11111110, 
    8'b00001111, 8'b10000000, 8'b00000001, 8'b11100000, 
    8'b00011111, 8'b10000000, 8'b00000001, 8'b11100000, 
    8'b00111111, 8'b10000000, 8'b00000001, 8'b11100000, 
    8'b01111111, 8'b10011111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b10011111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b10011111, 8'b11111111, 8'b11111110, 
    8'b01110111, 8'b10000011, 8'b10000001, 8'b11100000, 
    8'b00000111, 8'b10000111, 8'b11000001, 8'b11100000, 
    8'b00000111, 8'b10000111, 8'b11000001, 8'b11100000, 
    8'b00000111, 8'b10000011, 8'b11100001, 8'b11100000, 
    8'b00000111, 8'b10000001, 8'b11110001, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b11110001, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b01110001, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b00000001, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b00111111, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b00111111, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b00111111, 8'b11000000, 
    8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000
};

parameter [0:1023] char_ding={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00111100, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00111100, 
    8'b00111101, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11000000, 
    8'b00000011, 8'b11111111, 8'b11111111, 8'b11000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000001, 8'b10000011, 8'b11000000, 8'b00000000, 
    8'b00000001, 8'b11000011, 8'b11000000, 8'b00000000, 
    8'b00000011, 8'b11000011, 8'b11000000, 8'b00000000, 
    8'b00000011, 8'b11000011, 8'b11111111, 8'b11110000, 
    8'b00000011, 8'b11000011, 8'b11111111, 8'b11110000, 
    8'b00000111, 8'b11000011, 8'b11111111, 8'b11110000, 
    8'b00000111, 8'b10000011, 8'b11111111, 8'b11110000, 
    8'b00000111, 8'b11000011, 8'b11000000, 8'b00000000, 
    8'b00001111, 8'b11100011, 8'b11000000, 8'b00000000, 
    8'b00001111, 8'b11110011, 8'b11000000, 8'b00000000, 
    8'b00011111, 8'b11111011, 8'b11000000, 8'b00000000, 
    8'b00111110, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b01111110, 8'b01111111, 8'b11111100, 8'b00000110, 
    8'b01111100, 8'b00011111, 8'b11111111, 8'b11111110, 
    8'b01111000, 8'b00000111, 8'b11111111, 8'b11111110, 
    8'b01110000, 8'b00000000, 8'b01111111, 8'b11111110, 
    8'b00110000, 8'b00000000, 8'b00000000, 8'b00000000
};

parameter [0:1023] char_mo={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b10000001, 8'b11100011, 8'b11000000, 
    8'b00000111, 8'b10000001, 8'b11100011, 8'b11000000, 
    8'b00000111, 8'b10000001, 8'b11100011, 8'b11000000, 
    8'b00000111, 8'b10111111, 8'b11111111, 8'b11111110, 
    8'b00000111, 8'b10111111, 8'b11111111, 8'b11111110, 
    8'b00000111, 8'b10111111, 8'b11111111, 8'b11111110, 
    8'b00111111, 8'b11110001, 8'b11100011, 8'b11000000, 
    8'b01111111, 8'b11110001, 8'b11100011, 8'b11000000, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00000111, 8'b10001111, 8'b11111111, 8'b11111000, 
    8'b00001111, 8'b10001111, 8'b00000000, 8'b01111000, 
    8'b00001111, 8'b11001111, 8'b11111111, 8'b11111000, 
    8'b00001111, 8'b11101111, 8'b11111111, 8'b11111000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00011111, 8'b11111111, 8'b00000000, 8'b01111000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b01111111, 8'b10111111, 8'b11111111, 8'b11111000, 
    8'b11111111, 8'b10000000, 8'b00011100, 8'b00000000, 
    8'b01110111, 8'b10111111, 8'b11111111, 8'b11111110, 
    8'b01100111, 8'b10111111, 8'b11111111, 8'b11111110, 
    8'b01100111, 8'b10111111, 8'b11111111, 8'b11111110, 
    8'b00000111, 8'b10111111, 8'b11111111, 8'b11111110, 
    8'b00000111, 8'b10000001, 8'b11111111, 8'b10000000, 
    8'b00000111, 8'b10000011, 8'b11110111, 8'b11100000, 
    8'b00000111, 8'b10001111, 8'b11100011, 8'b11111000, 
    8'b00000111, 8'b10111111, 8'b11000001, 8'b11111110, 
    8'b00000111, 8'b10111111, 8'b10000000, 8'b11111110, 
    8'b00000111, 8'b10111100, 8'b00000000, 8'b00111110, 
    8'b00000011, 8'b10110000, 8'b00000000, 8'b00001100
};

parameter [0:1023] char_shi={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b01111000, 8'b11000000, 
    8'b00000000, 8'b00000000, 8'b01111011, 8'b11000000, 
    8'b00000000, 8'b00000000, 8'b01111011, 8'b11100000, 
    8'b00000000, 8'b00000000, 8'b01111001, 8'b11110000, 
    8'b00000000, 8'b00000000, 8'b01111000, 8'b11110000, 
    8'b00000000, 8'b00000000, 8'b01111000, 8'b11110000, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00111000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10111100, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10111100, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10111100, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10111100, 8'b00000000, 
    8'b00000000, 8'b11100000, 8'b00111100, 8'b00000000, 
    8'b00000000, 8'b11100000, 8'b00111110, 8'b00000000, 
    8'b00000000, 8'b11100000, 8'b00011110, 8'b00000000, 
    8'b00000000, 8'b11100000, 8'b00011110, 8'b00000000, 
    8'b00000000, 8'b11100000, 8'b00011110, 8'b00001000, 
    8'b00000000, 8'b11100000, 8'b11001111, 8'b00011110, 
    8'b00000000, 8'b11111111, 8'b11001111, 8'b00011110, 
    8'b00000111, 8'b11111111, 8'b11001111, 8'b10011110, 
    8'b01111111, 8'b11111111, 8'b11000111, 8'b10011110, 
    8'b01111111, 8'b11111110, 8'b00000111, 8'b11111100, 
    8'b00111111, 8'b10000000, 8'b00000011, 8'b11111100, 
    8'b00110000, 8'b00000000, 8'b00000001, 8'b11111000, 
    8'b00000000, 8'b00000000, 8'b00000001, 8'b11111000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00100000
};
parameter [0:1023] char_ji={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001100, 8'b00000000, 8'b00011110, 8'b00000000, 
    8'b00011110, 8'b00000000, 8'b00011110, 8'b00000000, 
    8'b00011111, 8'b00000000, 8'b00011110, 8'b00000000, 
    8'b00011111, 8'b11000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b11100000, 8'b00011110, 8'b00000000, 
    8'b00000011, 8'b11100000, 8'b00011110, 8'b00000000, 
    8'b00000001, 8'b11100000, 8'b00011110, 8'b00000000, 
    8'b00000000, 8'b11000000, 8'b00011110, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00011110, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00011110, 8'b00000000, 
    8'b01111111, 8'b10011111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b10011111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b10011111, 8'b11111111, 8'b11111110, 
    8'b00000111, 8'b10000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b10011000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b11111000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b11111000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b11111000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b11110000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b11100000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b00000000, 8'b00011110, 8'b00000000, 
    8'b00000010, 8'b00000000, 8'b00011110, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00011110, 8'b00000000
};
parameter [0:1023] char_suan={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00111100, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00111100, 8'b00000000, 
    8'b00001111, 8'b11111111, 8'b01111111, 8'b11111110, 
    8'b00001111, 8'b11111111, 8'b01111111, 8'b11111110, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00111110, 8'b01111001, 8'b11110011, 8'b11000000, 
    8'b01111100, 8'b01111001, 8'b11110011, 8'b11100000, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b00000000, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b00000000, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000000, 8'b01111000, 8'b00001111, 8'b00000000, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00000001, 8'b11110000, 8'b00001111, 8'b00000000, 
    8'b00000011, 8'b11110000, 8'b00001111, 8'b00000000, 
    8'b00011111, 8'b11100000, 8'b00001111, 8'b00000000, 
    8'b00011111, 8'b11000000, 8'b00001111, 8'b00000000, 
    8'b00001111, 8'b00000000, 8'b00001111, 8'b00000000, 
    8'b00001100, 8'b00000000, 8'b00001110, 8'b00000000
};
parameter [0:1023] char_xue={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b00000111, 8'b00000001, 8'b11100000, 
    8'b00001111, 8'b00001111, 8'b00000001, 8'b11100000, 
    8'b00001111, 8'b10001111, 8'b10000011, 8'b11100000, 
    8'b00000111, 8'b11000111, 8'b11000011, 8'b11100000, 
    8'b00000011, 8'b11000011, 8'b11000111, 8'b11000000, 
    8'b00000011, 8'b11100011, 8'b11000111, 8'b11000000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111000, 8'b00000000, 8'b00000000, 8'b00011100, 
    8'b00111001, 8'b11111111, 8'b11111111, 8'b10011100, 
    8'b00111001, 8'b11111111, 8'b11111111, 8'b10011100, 
    8'b00111001, 8'b11111111, 8'b11111111, 8'b10011100, 
    8'b00111001, 8'b11111111, 8'b11111111, 8'b10011100, 
    8'b00000000, 8'b00000000, 8'b01111111, 8'b00000000, 
    8'b00000000, 8'b00000001, 8'b11111100, 8'b00000000, 
    8'b00000000, 8'b00000001, 8'b11111000, 8'b00000000, 
    8'b00000000, 8'b00000001, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00000000, 8'b00000001, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000001, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000001, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00111111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00111111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00111111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00111111, 8'b00000000, 8'b00000000
};
parameter [0:1023] char_xi={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11110000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11110000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11110000, 
    8'b00001111, 8'b11111111, 8'b11111111, 8'b11110000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b11110000, 
    8'b00000001, 8'b10000000, 8'b00000000, 8'b11110000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b11110000, 
    8'b00000111, 8'b11100000, 8'b00000000, 8'b11110000, 
    8'b00000011, 8'b11110000, 8'b00000000, 8'b11110000, 
    8'b00000001, 8'b11111000, 8'b00000000, 8'b11110000, 
    8'b00000000, 8'b11111100, 8'b00000000, 8'b11110000, 
    8'b00000000, 8'b00111110, 8'b00000000, 8'b11110000, 
    8'b00000000, 8'b00011110, 8'b00000000, 8'b11110000, 
    8'b00000000, 8'b00001100, 8'b00011000, 8'b11110000, 
    8'b00000000, 8'b00000000, 8'b01111100, 8'b11110000, 
    8'b00000000, 8'b00000001, 8'b11111100, 8'b11110000, 
    8'b00000000, 8'b00000111, 8'b11111100, 8'b11110000, 
    8'b00000000, 8'b00011111, 8'b11110000, 8'b11110000, 
    8'b00000000, 8'b11111111, 8'b11000000, 8'b11110000, 
    8'b00000111, 8'b11111111, 8'b00000000, 8'b11110000, 
    8'b00011111, 8'b11111100, 8'b00000000, 8'b11110000, 
    8'b00011111, 8'b11100000, 8'b00000000, 8'b11100000, 
    8'b00011111, 8'b10000000, 8'b00000000, 8'b11100000, 
    8'b00011100, 8'b00000000, 8'b00000001, 8'b11100000, 
    8'b00000000, 8'b00000000, 8'b00000001, 8'b11100000, 
    8'b00000000, 8'b00000000, 8'b11111111, 8'b11100000, 
    8'b00000000, 8'b00000000, 8'b11111111, 8'b11000000, 
    8'b00000000, 8'b00000000, 8'b11111111, 8'b11000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};
parameter [0:1023] char_jing={
     8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00000000, 8'b11111000, 8'b00011111, 8'b00000000, 
    8'b00000000, 8'b01111000, 8'b00011110, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b00000001, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b00000001, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b00000001, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000011, 8'b11111111, 8'b11111111, 8'b11101000, 
    8'b00000000, 8'b00111110, 8'b01111000, 8'b00011110, 
    8'b00000000, 8'b01111100, 8'b01111000, 8'b00011110, 
    8'b00000000, 8'b11111100, 8'b01111000, 8'b00011110, 
    8'b00000111, 8'b11111000, 8'b01111100, 8'b00111110, 
    8'b01111111, 8'b11110000, 8'b00111111, 8'b11111110, 
    8'b01111111, 8'b11000000, 8'b00111111, 8'b11111100, 
    8'b01111111, 8'b00000000, 8'b00011111, 8'b11111000, 
    8'b00111000, 8'b00000000, 8'b00000000, 8'b00000000
};

parameter [0:1023] char_sai={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111100, 8'b00111100, 8'b00111000, 8'b00111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00000011, 8'b11111111, 8'b11111111, 8'b11000000, 
    8'b00000011, 8'b11111111, 8'b11111111, 8'b11000000, 
    8'b00000011, 8'b11111111, 8'b11111111, 8'b11000000, 
    8'b00000011, 8'b11111111, 8'b11111111, 8'b11000000, 
    8'b00000000, 8'b00111100, 8'b00111000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00000011, 8'b11110000, 8'b00001111, 8'b11000000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00111001, 8'b11000011, 8'b11000011, 8'b10011100, 
    8'b00000001, 8'b11000011, 8'b11000011, 8'b10000000, 
    8'b00000001, 8'b11000011, 8'b10000011, 8'b10000000, 
    8'b00000001, 8'b11000111, 8'b10000011, 8'b10000000, 
    8'b00000001, 8'b11000111, 8'b11110011, 8'b10000000, 
    8'b00000001, 8'b11001111, 8'b11111111, 8'b10000000, 
    8'b00000000, 8'b00111111, 8'b11111111, 8'b11000000, 
    8'b00001111, 8'b11111111, 8'b00111111, 8'b11110000, 
    8'b00011111, 8'b11111100, 8'b00000111, 8'b11110000, 
    8'b00001111, 8'b11111000, 8'b00000001, 8'b11110000, 
    8'b00001111, 8'b00000000, 8'b00000000, 8'b01100000
};

parameter [0:1023] char_yan={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b01111110, 8'b00111111, 8'b11111111, 8'b11111110, 
    8'b00111111, 8'b00111111, 8'b11111111, 8'b11111110, 
    8'b00011111, 8'b10111111, 8'b11111111, 8'b11111110, 
    8'b00001111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00000111, 8'b11111000, 8'b00000000, 8'b00011110, 
    8'b00000011, 8'b10111111, 8'b11111111, 8'b11111110, 
    8'b00110000, 8'b00111111, 8'b11111111, 8'b11111110, 
    8'b01111000, 8'b00111111, 8'b11111111, 8'b11111100, 
    8'b01111110, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b01111111, 8'b00011111, 8'b11111111, 8'b11111000, 
    8'b00011111, 8'b10011111, 8'b11111111, 8'b11111000, 
    8'b00001111, 8'b10011111, 8'b11111111, 8'b11111000, 
    8'b00000111, 8'b10011111, 8'b11111111, 8'b11111000, 
    8'b00000011, 8'b00011110, 8'b00111100, 8'b00111000, 
    8'b00000000, 8'b00011111, 8'b11111111, 8'b11111000, 
    8'b00000011, 8'b10011111, 8'b11111111, 8'b11111000, 
    8'b00000011, 8'b11011111, 8'b11111111, 8'b11111000, 
    8'b00000111, 8'b11011110, 8'b00111100, 8'b00111000, 
    8'b00000111, 8'b10011110, 8'b00111100, 8'b00111000, 
    8'b00000111, 8'b10011111, 8'b11111111, 8'b11111000, 
    8'b00001111, 8'b00011111, 8'b11111111, 8'b11111000, 
    8'b00001111, 8'b00011111, 8'b11111111, 8'b11111000, 
    8'b00011110, 8'b00000001, 8'b11000011, 8'b10000000, 
    8'b00011110, 8'b00000111, 8'b11100011, 8'b11100000, 
    8'b00111100, 8'b00011111, 8'b11100011, 8'b11111000, 
    8'b00111100, 8'b01111111, 8'b10000001, 8'b11111110, 
    8'b01111100, 8'b11111111, 8'b00000000, 8'b01111111, 
    8'b00111000, 8'b01111100, 8'b00000000, 8'b00011110, 
    8'b00000000, 8'b00110000, 8'b00000000, 8'b00000100
};
parameter [0:1023] char_shi2={
     8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000001, 8'b10000000, 
    8'b00000011, 8'b11000011, 8'b11000111, 8'b10000000, 
    8'b00000011, 8'b11000011, 8'b11000011, 8'b11000000, 
    8'b00000011, 8'b11000011, 8'b11000011, 8'b11100000, 
    8'b00000111, 8'b10000011, 8'b11000001, 8'b11100000, 
    8'b00000111, 8'b10000011, 8'b11000001, 8'b11110000, 
    8'b00001111, 8'b10000011, 8'b11000000, 8'b11110000, 
    8'b00001111, 8'b00000011, 8'b11000000, 8'b11111000, 
    8'b00011111, 8'b00000011, 8'b11000000, 8'b01111000, 
    8'b00111110, 8'b00000011, 8'b11000000, 8'b01111100, 
    8'b00111110, 8'b00000011, 8'b11000000, 8'b00111100, 
    8'b01111100, 8'b00000011, 8'b11000000, 8'b00111110, 
    8'b01111000, 8'b01111111, 8'b11000000, 8'b00011110, 
    8'b00011000, 8'b01111111, 8'b11000000, 8'b00011000, 
    8'b00000000, 8'b01111111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};
parameter [0:1023] char_dui={
     8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b11110000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b11110000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b11110000, 
    8'b00111111, 8'b11111100, 8'b00000000, 8'b11110000, 
    8'b00111111, 8'b11111100, 8'b00000000, 8'b11110000, 
    8'b00111111, 8'b11111100, 8'b00000000, 8'b11110000, 
    8'b00111111, 8'b11111101, 8'b11111111, 8'b11111110, 
    8'b00000000, 8'b00011101, 8'b11111111, 8'b11111110, 
    8'b00011000, 8'b00111101, 8'b11111111, 8'b11111110, 
    8'b00111000, 8'b00111101, 8'b11111111, 8'b11111110, 
    8'b00111100, 8'b00111100, 8'b00000000, 8'b11110000, 
    8'b00111110, 8'b00111100, 8'b00000000, 8'b11110000, 
    8'b00011111, 8'b00111000, 8'b11000000, 8'b11110000, 
    8'b00001111, 8'b11111001, 8'b11100000, 8'b11110000, 
    8'b00001111, 8'b11111001, 8'b11100000, 8'b11110000, 
    8'b00000111, 8'b11110001, 8'b11110000, 8'b11110000, 
    8'b00000011, 8'b11110000, 8'b11111000, 8'b11110000, 
    8'b00000001, 8'b11110000, 8'b01111000, 8'b11110000, 
    8'b00000001, 8'b11111000, 8'b01111100, 8'b11110000, 
    8'b00000011, 8'b11111000, 8'b00111110, 8'b11110000, 
    8'b00000111, 8'b11111100, 8'b00011110, 8'b11110000, 
    8'b00000111, 8'b11111110, 8'b00011000, 8'b11110000, 
    8'b00001111, 8'b10011110, 8'b00000000, 8'b11110000, 
    8'b00011111, 8'b00011110, 8'b00000000, 8'b11110000, 
    8'b00111110, 8'b00001100, 8'b00000000, 8'b11110000, 
    8'b01111100, 8'b00000000, 8'b00000000, 8'b11110000, 
    8'b01111000, 8'b00000000, 8'b00000000, 8'b11110000, 
    8'b01110000, 8'b00000000, 8'b01111111, 8'b11100000, 
    8'b00100000, 8'b00000000, 8'b01111111, 8'b11100000, 
    8'b00000000, 8'b00000000, 8'b00111111, 8'b11100000, 
    8'b00000000, 8'b00000000, 8'b00111111, 8'b10000000
};

parameter [0:1023] char_cuo={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b00000000, 8'b01110000, 8'b11100000, 
    8'b00001111, 8'b00000000, 8'b01110000, 8'b11100000, 
    8'b00001111, 8'b00000000, 8'b01110000, 8'b11100000, 
    8'b00001111, 8'b00000000, 8'b01110000, 8'b11100000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00111100, 8'b00000000, 8'b01110000, 8'b11100000, 
    8'b00111100, 8'b00000000, 8'b01110000, 8'b11100000, 
    8'b01111000, 8'b00000000, 8'b01110000, 8'b11100000, 
    8'b11111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b11111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00001111, 8'b11110000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000001, 8'b11111111, 8'b11111000, 
    8'b00000011, 8'b11000001, 8'b11111111, 8'b11111000, 
    8'b00111111, 8'b11111101, 8'b11111111, 8'b11111000, 
    8'b00111111, 8'b11111101, 8'b11111111, 8'b11111000, 
    8'b00111111, 8'b11111101, 8'b11000000, 8'b00111000, 
    8'b00111111, 8'b11111101, 8'b11000000, 8'b00111000, 
    8'b00000011, 8'b11000001, 8'b11111111, 8'b11111000, 
    8'b00000011, 8'b11000001, 8'b11111111, 8'b11111000, 
    8'b00000011, 8'b11000001, 8'b11111111, 8'b11111000, 
    8'b00000011, 8'b11000001, 8'b11000000, 8'b00111000, 
    8'b00000011, 8'b11011101, 8'b11000000, 8'b00111000, 
    8'b00000011, 8'b11111111, 8'b11000000, 8'b00111000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00000111, 8'b11111001, 8'b11111111, 8'b11111000, 
    8'b00000111, 8'b11100001, 8'b11111111, 8'b11111000, 
    8'b00000011, 8'b00000001, 8'b11000000, 8'b00111000, 
    8'b00000000, 8'b00000001, 8'b11000000, 8'b00111000
};*/

    wire [9:0] pix_x;
    wire [9:0] pix_y;
    wire vga_clk; //25MHz
    wire [15:0] pix_data;
    wire rst_n;
    assign rst_n= reset_n;
    assign vga_clk = clk;
    /*clk_wiz_0 clk_inst(   // clk_wiz_0 used ip core
        .clk_in1(clk),
        .reset(~rst_n),
        .clk_out1(vga_clk)
    );*/

    // horizontal counter
    reg [9:0] hc;
    always @(posedge vga_clk) begin
        if (~rst_n) hc <= 0;
        else if (hc == `H_LINE_PERIOD - 1) hc <= 0;
        else hc <= hc + 1;
    end

    // vertical counter
    reg [9:0] vc;
    always @(posedge vga_clk) begin
        if (~rst_n) vc <= 0;
        else if (vc == `V_FRAME_PERIOD - 1) vc <= 0;
        else if (hc == `H_LINE_PERIOD - 1) vc <= vc + 1;
        else vc <= vc;
    end

    wire [9:0] hc0, vc0;
    assign hsync = (hc < `H_SYNC_PULSE) ? 0 : 1;
    assign vsync = (vc < `V_SYNC_PULSE) ? 0 : 1;
    assign hc0 = hc - `H_SYNC_PULSE - `H_BACK_PORCH;
    assign vc0 = vc - `V_SYNC_PULSE - `V_BACK_PORCH;

    wire active;  // is the point active
    assign active = (hc >= `H_SYNC_PULSE + `H_BACK_PORCH) &&
                    (hc < `H_SYNC_PULSE + `H_BACK_PORCH + `H_ACTIVE_TIME) &&
                    (vc >= `V_SYNC_PULSE + `V_BACK_PORCH) &&
                    (vc < `V_SYNC_PULSE + `V_BACK_PORCH + `V_ACTIVE_TIME) ? 1 : 0;

    reg [10:0] idx;
    
    ///bcd///
   /* wire [0:1023]  bcd_0;
    wire [0:1023]  bcd_1;
    wire [0:1023]  bcd_2;
    wire [0:1023]  bcd_3;
    wire [0:1023]  bcd_4;
    wire [0:1023]  bcd_5;
    wire [0:1023]  bcd_6;
    wire [0:1023]  bcd_7;*/
    /*vga_decoder_8 vga_decoder_8_inst_0(
        .seg(segment0),
        .vga(bcd_0)
    );
    vga_decoder_8 vga_decoder_8_inst_1(
        .seg(segment1),
        .vga(bcd_1)
    );
    vga_decoder_8 vga_decoder_8_inst_2(
        .seg(segment2),
        .vga(bcd_2)
    );
    vga_decoder_8 vga_decoder_8_inst_3(
        .seg(segment3),
        .vga(bcd_3)
    );
    vga_decoder_8 vga_decoder_8_inst_4(
        .seg(segment4),
        .vga(bcd_4)
    );
    vga_decoder_8 vga_decoder_8_inst_5(
        .seg(segment5),
        .vga(bcd_5)
    );
    vga_decoder_8 vga_decoder_8_inst_6(
        .seg(segment6),
        .vga(bcd_6)
    );
    vga_decoder_8 vga_decoder_8_inst_7(
        .seg(segment7),
        .vga(bcd_7)
    );*/
    


    always @(*) begin
        if (~rst_n) begin
            red = 0;
            green = 0;
            blue = 0;
        end
        else if (active) begin
            ///game_mode///
            if (hc0 >= 480 + 0*`char_width && hc0 < 480 + 1*`char_width && vc0 >= 32 && vc0 < 32 + `char_width) begin
                idx = hc0 - 480 + 32 * (vc0 - 32);
                /*if (game_mode ==`power_off) begin
                    if (char_guan[idx] == 1) {red, green, blue} = `WHITE;
                    else {red, green, blue} = `BLACK;
                end
                else if (game_mode ==`stand_by) begin
                    if (char_dai[idx] == 1) {red, green, blue} = `WHITE;
                    else {red, green, blue} = `BLACK;
                end
                // else if (game_mode ==`idle) begin
                //     if (char_zou[idx] == 1) {red, green, blue} = `WHITE;
                //     else {red, green, blue} = `BLACK;
                // end
                else if (game_mode ==`calc_mode) begin
                    if (char_ji[idx] == 1) {red, green, blue} = `WHITE;
                    else {red, green, blue} = `BLACK;
                end
                else if (game_mode ==`learn_mode) begin
                    if (char_xue[idx] == 1) {red, green, blue} = `WHITE;
                    else {red, green, blue} = `BLACK;
                end
                else if (game_mode ==`competition_mode) begin
                    if (char_jing[idx] == 1) {red, green, blue} = `WHITE;
                    else {red, green, blue} = `BLACK;
                end
                else if (game_mode ==`demonstration_mode) begin
                    if (char_yan[idx] == 1) {red, green, blue} = `WHITE;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    {red, green, blue} = `BLACK;
                end
                
            end
            else if (hc0 >= 480 + 1*`char_width && hc0 < 480 + 2*`char_width && vc0 >= 32 && vc0 < 32 + `char_width) begin
                idx = hc0 - 480 -`char_width + 32 * (vc0 - 32);
                if (game_mode ==`power_off) begin
                    if (char_ji2[idx] == 1) {red, green, blue} = `WHITE;
                    else {red, green, blue} = `BLACK;
                end
                else if (game_mode ==`stand_by) begin
                    if (char_ding[idx] == 1) {red, green, blue} = `WHITE;
                    else {red, green, blue} = `BLACK;
                end
                else if (game_mode==`calc_mode) begin
                    if(char_suan[idx] == 1) {red, green, blue} = `WHITE;
                    else {red, green, blue} = `BLACK;
                end
                else if (game_mode==`learn_mode) begin
                    if(char_xi[idx] == 1) {red, green, blue} = `WHITE;
                    else {red, green, blue} = `BLACK;
                end
                else if (game_mode==`competition_mode) begin
                    if(char_sai[idx] == 1) {red, green, blue} = `WHITE;
                    else {red, green, blue} = `BLACK;
                end
                else if (game_mode==`demonstration_mode) begin
                    if(char_shi2[idx] == 1) {red, green, blue} = `WHITE;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    {red, green, blue} = `BLACK;
                end*/
                
            end
            /*else if (hc0 >= 480 + 2*`char_width && hc0 < 480 + 3*`char_width && vc0 >= 32 && vc0 < 32 + `char_width) begin
                /*idx = hc0 - 480 - 2*`char_width + 32 * (vc0 - 32);
                if (char_mo[idx] == 1) {red, green, blue} = `WHITE;
                else {red, green, blue} = `BLACK;
            end*/
            else if (hc0 >= 480 + 3*`char_width && hc0 < 480 + 4*`char_width && vc0 >= 32 && vc0 < 32 + `char_width) begin
                /*idx = hc0 - 480 - 3*`char_width + 32 * (vc0 - 32);
                if (char_shi[idx] == 1) {red, green, blue} = `WHITE;
                else {red, green, blue} = `BLACK;*/
            end
            ///switches///
            else if (hc0 >= 96 + 0*`char_width && hc0<96 + 1*`char_width && vc0 >= 128 && vc0 < 128 + `char_width) begin
                idx = hc0 - 96 + 32 * (vc0 - 128);
                /*if (script[7] == 1) begin
                    if (num_one[idx]){red, green, blue} = `RED;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `RED;
                    else {red, green, blue} = `BLACK;
                end*/
            end
            else if (hc0 >= 96 + 1*`char_width && hc0<96 + 2*`char_width && vc0 >= 128 && vc0 < 128 + `char_width) begin
                idx = hc0 - 96 - `char_width + 32 * (vc0 - 128);
                /*if (script[6] == 1) begin
                    if (num_one[idx]){red, green, blue} = `RED;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `RED;
                    else {red, green, blue} = `BLACK;
                end*/
            end
            else if (hc0 >= 96 + 2*`char_width && hc0<96 + 3*`char_width && vc0 >= 128 && vc0 < 128 + `char_width) begin
                idx = hc0 - 96 - 2*`char_width + 32 * (vc0 - 128);
                /*if (script[5] == 1) begin
                    if (num_one[idx]){red, green, blue} = `RED;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `RED;
                    else {red, green, blue} = `BLACK;
                end*/
            end
            else if (hc0 >= 96 + 3*`char_width && hc0<96 + 4*`char_width && vc0 >= 128 && vc0 < 128 + `char_width) begin
                idx = hc0 - 96 - 3*`char_width + 32 * (vc0 - 128);
                /*if (script[4] == 1) begin
                    if (num_one[idx]){red, green, blue} = `RED;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `RED;
                    else {red, green, blue} = `BLACK;
                end*/
            end
            else if (hc0 >= 96 + 4*`char_width && hc0<96 + 5*`char_width && vc0 >= 128 && vc0 < 128 + `char_width) begin
                idx = hc0 - 96 - 4*`char_width + 32 * (vc0 - 128);
                /*if (script[3] == 1) begin
                    if (num_one[idx]){red, green, blue} = `RED;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `RED;
                    else {red, green, blue} = `BLACK;
                end*/
            end
            else if (hc0 >= 96 + 5*`char_width && hc0<96 + 6*`char_width && vc0 >= 128 && vc0 < 128 + `char_width) begin
                idx = hc0 - 96 - 5*`char_width + 32 * (vc0 - 128);
                /*if (script[2] == 1) begin
                    if (num_one[idx]){red, green, blue} = `RED;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `RED;
                    else {red, green, blue} = `BLACK;
                end
            end
            else if (hc0 >= 96 + 6*`char_width && hc0<96 + 7*`char_width && vc0 >= 128 && vc0 < 128 + `char_width) begin
                idx = hc0 - 96 - 6*`char_width + 32 * (vc0 - 128);
                if (script[1] == 1) begin
                    if (num_one[idx]){red, green, blue} = `RED;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `RED;
                    else {red, green, blue} = `BLACK;
                end
            end
            else if (hc0 >= 96 + 7*`char_width && hc0<96 + 8*`char_width && vc0 >= 128 && vc0 < 128 + `char_width) begin
                idx = hc0 - 96 - 7*`char_width + 32 * (vc0 - 128);
                if (script[0] == 1) begin
                    if (num_one[idx]){red, green, blue} = `RED;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `RED;
                    else {red, green, blue} = `BLACK;
                end
            end*/
            end
            ///led_1///
            else if (hc0 >= 96 + 0*`char_width && hc0<96 + 1*`char_width && vc0 >= 256 && vc0 < 256 + `char_width) begin
                idx = hc0 - 96 + 32 * (vc0 - 256);
                if (data[7] == 1) begin
                    if (num_one[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
            end
            else if (hc0 >= 96 + 1*`char_width && hc0<96 + 2*`char_width && vc0 >= 256 && vc0 < 256 + `char_width) begin
                idx = hc0 - 96 - `char_width + 32 * (vc0 - 256);
                if (data[6] == 1) begin
                    if (num_one[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
            end
            else if (hc0 >= 96 + 2*`char_width && hc0<96 + 3*`char_width && vc0 >= 256 && vc0 < 256 + `char_width) begin
                idx = hc0 - 96 - 2*`char_width + 32 * (vc0 - 256);
                if (data[5] == 1) begin
                    if (num_one[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
            end
            else if (hc0 >= 96 + 3*`char_width && hc0<96 + 4*`char_width && vc0 >= 256 && vc0 < 256 + `char_width) begin
                idx = hc0 - 96 - 3*`char_width + 32 * (vc0 - 256);
                if (data[4] == 1) begin
                    if (num_one[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
            end
            else if (hc0 >= 96 + 4*`char_width && hc0<96 + 5*`char_width && vc0 >= 256 && vc0 < 256 + `char_width) begin
                idx = hc0 - 96 - 4*`char_width + 32 * (vc0 - 256);
                if (data[3] == 1) begin
                    if (num_one[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
            end
            else if (hc0 >= 96 + 5*`char_width && hc0<96 + 6*`char_width && vc0 >= 256 && vc0 < 256 + `char_width) begin
                idx = hc0 - 96 - 5*`char_width + 32 * (vc0 - 256);
                if (data[2] == 1) begin
                    if (num_one[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
            end
            else if (hc0 >= 96 + 6*`char_width && hc0<96 + 7*`char_width && vc0 >= 256 && vc0 < 256 + `char_width) begin
                idx = hc0 - 96 - 6*`char_width + 32 * (vc0 - 256);
                if (data[1] == 1) begin
                    if (num_one[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
            end
            else if (hc0 >= 96 + 7*`char_width && hc0<96 + 8*`char_width && vc0 >= 256 && vc0 < 256 + `char_width) begin
                idx = hc0 - 96 - 7*`char_width + 32 * (vc0 - 256);
                if (data[0] == 1) begin
                    if (num_one[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
            end
            ///led_2///
            /*
            else if (hc0 >= 96 + 0*`char_width && hc0<96 + 1*`char_width && vc0 >= 320 && vc0 < 320 + `char_width) begin
                idx = hc0 - 96 + 32 * (vc0 - 320);
                if (led_2[7] == 1) begin
                    if (num_one[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
            end
            else if (hc0 >= 96 + 1*`char_width && hc0<96 + 2*`char_width && vc0 >= 320 && vc0 < 320 + `char_width) begin
                idx = hc0 - 96 - `char_width + 32 * (vc0 - 320);
                if (led_2[6] == 1) begin
                    if (num_one[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
            end
            else if (hc0 >= 96 + 2*`char_width && hc0<96 + 3*`char_width && vc0 >= 320 && vc0 < 320 + `char_width) begin
                idx = hc0 - 96 - 2*`char_width + 32 * (vc0 - 320);
                if (led_2[5] == 1) begin
                    if (num_one[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
            end
            else if (hc0 >= 96 + 3*`char_width && hc0<96 + 4*`char_width && vc0 >= 320 && vc0 < 320 + `char_width) begin
                idx = hc0 - 96 - 3*`char_width + 32 * (vc0 - 320);
                if (led_2[4] == 1) begin
                    if (num_one[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
            end
            else if (hc0 >= 96 + 4*`char_width && hc0<96 + 5*`char_width && vc0 >= 320 && vc0 < 320 + `char_width) begin
                idx = hc0 - 96 - 4*`char_width + 32 * (vc0 - 320);
                if (led_2[3] == 1) begin
                    if (num_one[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
            end
            else if (hc0 >= 96 + 5*`char_width && hc0<96 + 6*`char_width && vc0 >= 320 && vc0 < 320 + `char_width) begin
                idx = hc0 - 96 - 5*`char_width + 32 * (vc0 - 320);
                if (led_2[2] == 1) begin
                    if (num_one[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
            end
            else if (hc0 >= 96 + 6*`char_width && hc0<96 + 7*`char_width && vc0 >= 320 && vc0 < 320 + `char_width) begin
                idx = hc0 - 96 - 6*`char_width + 32 * (vc0 - 320);
                if (led_2[1] == 1) begin
                    if (num_one[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
            end
            else if (hc0 >= 96 + 7*`char_width && hc0<96 + 8*`char_width && vc0 >= 320 && vc0 < 320 + `char_width) begin
                idx = hc0 - 96 - 7*`char_width + 32 * (vc0 - 320);
                if (led_2[0] == 1) begin
                    if (num_one[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
                else begin
                    if (num_zero[idx]){red, green, blue} = `GREEN;
                    else {red, green, blue} = `BLACK;
                end
            end
            ///BCD///
            else if (hc0 >= 96 + 0*`char_width && hc0<96 + 1*`char_width && vc0 >= 384 && vc0 < 384 + `char_width) begin
                idx = hc0 - 96 + 32 * (vc0 - 384);
                if (bcd_7[idx] == 1) {red, green, blue} = `GOLDEN;
                else {red, green, blue} = `BLACK;
            end
            else if (hc0 >= 96 + 1*`char_width && hc0<96 + 2*`char_width && vc0 >= 384 && vc0 < 384 + `char_width) begin
                idx = hc0 - 96 - `char_width + 32 * (vc0 - 384);
                if (bcd_6[idx] == 1) {red, green, blue} = `GOLDEN;
                else {red, green, blue} = `BLACK;
            end
            else if (hc0 >= 96 + 2*`char_width && hc0<96 + 3*`char_width && vc0 >= 384 && vc0 < 384 + `char_width) begin
                idx = hc0 - 96 - 2*`char_width + 32 * (vc0 - 384);
                if (bcd_5[idx] == 1) {red, green, blue} = `GOLDEN;
                else {red, green, blue} = `BLACK;
            end
            else if (hc0 >= 96 + 3*`char_width && hc0<96 + 4*`char_width && vc0 >= 384 && vc0 < 384 + `char_width) begin
                idx = hc0 - 96 - 3*`char_width + 32 * (vc0 - 384);
                if (bcd_4[idx] == 1) {red, green, blue} = `GOLDEN;
                else {red, green, blue} = `BLACK;
            end
            else if (hc0 >= 96 + 4*`char_width && hc0<96 + 5*`char_width && vc0 >= 384 && vc0 < 384 + `char_width) begin
                idx = hc0 - 96 - 4*`char_width + 32 * (vc0 - 384);
                if (bcd_3[idx] == 1) {red, green, blue} = `GOLDEN;
                else {red, green, blue} = `BLACK;
            end
            else if (hc0 >= 96 + 5*`char_width && hc0<96 + 6*`char_width && vc0 >= 384 && vc0 < 384 + `char_width) begin
                idx = hc0 - 96 - 5*`char_width + 32 * (vc0 - 384);
                if (bcd_2[idx] == 1) {red, green, blue} = `GOLDEN;
                else {red, green, blue} = `BLACK;
            end
            else if (hc0 >= 96 + 6*`char_width && hc0<96 + 7*`char_width && vc0 >= 384 && vc0 < 384 + `char_width) begin
                idx = hc0 - 96 - 6*`char_width + 32 * (vc0 - 384);
                if (bcd_1[idx] == 1) {red, green, blue} = `GOLDEN;
                else {red, green, blue} = `BLACK;
            end
            else if (hc0 >= 96 + 7*`char_width && hc0<96 + 8*`char_width && vc0 >= 384 && vc0 < 384 + `char_width) begin
                idx = hc0 - 96 - 7*`char_width + 32 * (vc0 - 384);
                if (bcd_0[idx] == 1) {red, green, blue} = `GOLDEN;
                else {red, green, blue} = `BLACK;
            end
            else begin
                {red, green, blue} = `BLACK;
            end
        end*/
        else begin
            {red, green, blue} = `BLACK;
        end
    end
end
            

endmodule