`timescale 1ns/1ps
`include "Constants.vh"

// Module: IF
// Description: Instruction Fetch stage. This module uses an ICache to get instructions and integrates
// the ImmGenerator and Branch_Predictor modules to update the Program Counter (PC)
// based on branch signals and predictions.
module IF (
    input         clk,         // Clock signal
    input         rst,         // Reset signal (active high)
    // Pipeline control:
    input         IF_ID_Write,   // Enable writing to IF/ID pipeline register
    input         Branch,      // External branch signal from EX stage
    // ICache interface:
    output [31:0] MemPC,       // Address passed to the ICache module
    input  [31:0] MemInst,     // Instruction returned from ICache
    output        ICacheStall, // Stall signal from ICache module
    // Outputs to the next pipeline stage:
    output reg [31:0] PcOut,   // PC passed to the IF/ID pipeline register
    output reg [31:0] InstOut  // Fetched instruction passed to the IF/ID pipeline register
);

  // Internal PC register used to track the current PC
  reg [31:0] PC;
  
  // Immediate value generated by ImmGenerator
  wire [31:0] Imm32;
  
  // Branch_Predictor module outputs
  wire        BpPredictFail;
  wire [31:0] BpTargetPC;
  wire        BpPredictResult;
  
  // Determine if the instruction is a jump or branch instruction
  wire Jump;
  wire BranchInst;
  wire Predict;
  assign Jump = ((MemInst[6:0] == `JAL_OPERATION) || (MemInst[6:0] == `JALR_OPERATION));
  assign BranchInst = ((MemInst[6:0] == `BRANCH_OPERATION) || Jump);
  // Use branch prediction only for conditional branches (non-jump)
  assign Predict = (~Jump) & BranchInst;
  
  // Instantiate the Branch_Predictor module
  Branch_Predictor BP (
      .clk(clk),
      .rst(rst),
      .stall(ICacheStall),
      .branch(BranchInst),
      .predict(Predict),
      .excp(1'b0),            // No exception handling in IF stage
      .sret(1'b0),
      // If jump, use 0 for rs1; otherwise use bits [19:15] of the instruction
      .rs1( Jump ? 5'd0 : MemInst[19:15]),
      .rd(MemInst[11:7]),
      .pc(PC),
      .imm(Imm32),
      // Use current PC as previous values in the update mechanism
      .old_pc(PC),
      .old_branch_pc(PC),
      .old_predict_pc(PC),
      .old_predict(1'b0),
      .old_actual(1'b0),
      .old_branch(1'b0),
      .target_pc(BpTargetPC),
      .predict_result(BpPredictResult),
      .predict_fail(BpPredictFail)
  );
  
  // Instantiate the ImmGenerator module
  ImmGenerator ImmGen (
      .Instruction(MemInst),
      .ImmData(Imm32)
  );
  
  // Compute the next PC value using combinational logic.
  // If branch prediction fails, use the correct target PC.
  // Otherwise, if an external Branch signal is high, use PC + Imm32.
  // Otherwise, increment PC by 4.
  wire [31:0] NextPC;
  assign NextPC = BpPredictFail ? BpTargetPC : (Branch ? (PC + Imm32) : (PC + 32'd4));

  // Use a single always block to:
  // - Latch current PC into PcOut (and capture MemInst into InstOut)
  // - Update the internal PC to NextPC
  always @(posedge clk or posedge rst) begin
      if (rst) begin
          PC     <= 32'd0;
          PcOut  <= 32'd0;
          InstOut<= 32'd0;
      end else if (IF_ID_Write) begin
          // Latch current PC and fetched instruction into the IF/ID pipeline registers
          PcOut  <= PC;
          InstOut<= MemInst;
          // Update PC for the next cycle
          PC     <= NextPC;
      end
  end
  
  // Instantiate the ICache module.
  ICache U_Cache (
      .clk(clk),
      .rst(rst),
      .Addr(PC),
      .Inst(MemInst),
      .ICacheStall(ICacheStall),
      .MemPc(MemPC)
  );

endmodule